module jesd204_phy #() ();
    pcs ()
endmodule